`ifndef DEFINES
`define DEFINES

// BIOS width

`define BIOS_AWIDTH  12
`define BIOS_DWIDTH  32

// REGFILE width

`define REG_AWIDTH  32
`define REG_DWIDTH  32



// IMEM width
`define IMEM_AWIDTH  14
`define IMEM_DWIDTH  32

// DMEM_width
`define DMEM_AWIDTH  32
`define DMEM_DWIDTH  32

`define ALUOP_RTYPE 3'b000
`define ALUOP_

`endif

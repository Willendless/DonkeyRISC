`include "../defines.vh"
`include "../Opcode.vh"

module id_top (
    input wire[`IMEM_DWIDTH] inst_i,

    // data from regfile
    input wire[`]

)



endmodule
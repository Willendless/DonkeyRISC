/**
* execution stage of DonkeyRISCV
*   @OUTPUT:
*   
* 
*
*/
`include "../defines.vh"

module ex (
    
);

endmodule // ex 
module branch_comp(
    input [2:0] branch_type,
    input [31:0] reg1,
    input [31:0] imm1
);

endmodule
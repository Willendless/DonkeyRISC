`ifndef DEFINES
`define DEFINES

// BIOS width

`define BIOS_AWIDTH  12
`define BIOS_DWIDTH  32

// REGFILE width

`define REG_AWIDTH  32
`define REG_DWIDTH  32



// IMEM width
`define IMEM_AWIDTH  14
`define IMEM_DWIDTH  32

// DMEM_width
`define DMEM_AWIDTH  32
`define DMEM_DWIDTH  32

`define ALUOP_RTYPE 2'b00
`define ALUOP_ISTYPE 2'b01
`define ALUOP_OTHER 2'b10

`endif
